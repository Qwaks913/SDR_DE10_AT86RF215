// soc_system.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk_clk,                    //                    clk.clk
		output wire        hps_0_h2f_reset_reset_n,    //        hps_0_h2f_reset.reset_n
		output wire        hps_0_spim0_f_txd,          //          hps_0_spim0_f.txd
		input  wire        hps_0_spim0_f_rxd,          //                       .rxd
		input  wire        hps_0_spim0_f_ss_in_n,      //                       .ss_in_n
		output wire        hps_0_spim0_f_ssi_oe_n,     //                       .ssi_oe_n
		output wire        hps_0_spim0_f_ss_0_n,       //                       .ss_0_n
		output wire        hps_0_spim0_f_ss_1_n,       //                       .ss_1_n
		output wire        hps_0_spim0_f_ss_2_n,       //                       .ss_2_n
		output wire        hps_0_spim0_f_ss_3_n,       //                       .ss_3_n
		output wire        hps_0_spim0_sclk_out_f_clk, // hps_0_spim0_sclk_out_f.clk
		input  wire        lvds_clk_input_clk,         //         lvds_clk_input.clk
		input  wire [31:0] lvds_iq_hps_in_new_signal,  //         lvds_iq_hps_in.new_signal
		output wire [14:0] memory_mem_a,               //                 memory.mem_a
		output wire [2:0]  memory_mem_ba,              //                       .mem_ba
		output wire        memory_mem_ck,              //                       .mem_ck
		output wire        memory_mem_ck_n,            //                       .mem_ck_n
		output wire        memory_mem_cke,             //                       .mem_cke
		output wire        memory_mem_cs_n,            //                       .mem_cs_n
		output wire        memory_mem_ras_n,           //                       .mem_ras_n
		output wire        memory_mem_cas_n,           //                       .mem_cas_n
		output wire        memory_mem_we_n,            //                       .mem_we_n
		output wire        memory_mem_reset_n,         //                       .mem_reset_n
		inout  wire [31:0] memory_mem_dq,              //                       .mem_dq
		inout  wire [3:0]  memory_mem_dqs,             //                       .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,           //                       .mem_dqs_n
		output wire        memory_mem_odt,             //                       .mem_odt
		output wire [3:0]  memory_mem_dm,              //                       .mem_dm
		input  wire        memory_oct_rzqin,           //                       .oct_rzqin
		input  wire        reset_reset_n,              //                  reset.reset_n
		input  wire        word_valid_word_valid       //             word_valid.word_valid
	);

	wire    [1:0] hps_0_h2f_axi_master_awburst;                            // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire    [3:0] hps_0_h2f_axi_master_arlen;                              // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire    [7:0] hps_0_h2f_axi_master_wstrb;                              // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_wready;                             // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [11:0] hps_0_h2f_axi_master_rid;                                // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_rready;                             // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire    [3:0] hps_0_h2f_axi_master_awlen;                              // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire   [11:0] hps_0_h2f_axi_master_wid;                                // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire    [3:0] hps_0_h2f_axi_master_arcache;                            // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire          hps_0_h2f_axi_master_wvalid;                             // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire   [29:0] hps_0_h2f_axi_master_araddr;                             // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire    [2:0] hps_0_h2f_axi_master_arprot;                             // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire    [2:0] hps_0_h2f_axi_master_awprot;                             // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire   [63:0] hps_0_h2f_axi_master_wdata;                              // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_arvalid;                            // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire    [3:0] hps_0_h2f_axi_master_awcache;                            // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire   [11:0] hps_0_h2f_axi_master_arid;                               // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire    [1:0] hps_0_h2f_axi_master_arlock;                             // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire    [1:0] hps_0_h2f_axi_master_awlock;                             // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                             // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire    [1:0] hps_0_h2f_axi_master_bresp;                              // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire          hps_0_h2f_axi_master_arready;                            // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire   [63:0] hps_0_h2f_axi_master_rdata;                              // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire          hps_0_h2f_axi_master_awready;                            // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                            // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire    [2:0] hps_0_h2f_axi_master_arsize;                             // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire          hps_0_h2f_axi_master_bready;                             // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire          hps_0_h2f_axi_master_rlast;                              // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire          hps_0_h2f_axi_master_wlast;                              // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire    [1:0] hps_0_h2f_axi_master_rresp;                              // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire   [11:0] hps_0_h2f_axi_master_awid;                               // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire   [11:0] hps_0_h2f_axi_master_bid;                                // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire          hps_0_h2f_axi_master_bvalid;                             // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire    [2:0] hps_0_h2f_axi_master_awsize;                             // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire          hps_0_h2f_axi_master_awvalid;                            // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire          hps_0_h2f_axi_master_rvalid;                             // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire   [63:0] mm_interconnect_0_mm_bridge_0_s0_readdata;               // mm_bridge_0:s0_readdata -> mm_interconnect_0:mm_bridge_0_s0_readdata
	wire          mm_interconnect_0_mm_bridge_0_s0_waitrequest;            // mm_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_bridge_0_s0_waitrequest
	wire          mm_interconnect_0_mm_bridge_0_s0_debugaccess;            // mm_interconnect_0:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	wire    [9:0] mm_interconnect_0_mm_bridge_0_s0_address;                // mm_interconnect_0:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	wire          mm_interconnect_0_mm_bridge_0_s0_read;                   // mm_interconnect_0:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	wire    [7:0] mm_interconnect_0_mm_bridge_0_s0_byteenable;             // mm_interconnect_0:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	wire          mm_interconnect_0_mm_bridge_0_s0_readdatavalid;          // mm_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_bridge_0_s0_readdatavalid
	wire          mm_interconnect_0_mm_bridge_0_s0_write;                  // mm_interconnect_0:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	wire   [63:0] mm_interconnect_0_mm_bridge_0_s0_writedata;              // mm_interconnect_0:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	wire    [0:0] mm_interconnect_0_mm_bridge_0_s0_burstcount;             // mm_interconnect_0:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                         // hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                           // hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                           // hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_wready;                          // mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                             // mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_rready;                          // hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                           // hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                             // hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                         // hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	wire          hps_0_h2f_lw_axi_master_wvalid;                          // hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                          // hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                          // hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                          // hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                           // hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_arvalid;                         // hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                         // hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                            // hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                          // hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                          // hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                          // hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                           // mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire          hps_0_h2f_lw_axi_master_arready;                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                           // mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire          hps_0_h2f_lw_axi_master_awready;                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                         // hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                          // hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	wire          hps_0_h2f_lw_axi_master_bready;                          // hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	wire          hps_0_h2f_lw_axi_master_rlast;                           // mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire          hps_0_h2f_lw_axi_master_wlast;                           // hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                           // mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                            // hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                             // mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire          hps_0_h2f_lw_axi_master_bvalid;                          // mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                          // hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	wire          hps_0_h2f_lw_axi_master_awvalid;                         // hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	wire          hps_0_h2f_lw_axi_master_rvalid;                          // mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire   [31:0] mm_interconnect_1_msgdma_0_csr_readdata;                 // msgdma_0:csr_readdata -> mm_interconnect_1:msgdma_0_csr_readdata
	wire    [2:0] mm_interconnect_1_msgdma_0_csr_address;                  // mm_interconnect_1:msgdma_0_csr_address -> msgdma_0:csr_address
	wire          mm_interconnect_1_msgdma_0_csr_read;                     // mm_interconnect_1:msgdma_0_csr_read -> msgdma_0:csr_read
	wire    [3:0] mm_interconnect_1_msgdma_0_csr_byteenable;               // mm_interconnect_1:msgdma_0_csr_byteenable -> msgdma_0:csr_byteenable
	wire          mm_interconnect_1_msgdma_0_csr_write;                    // mm_interconnect_1:msgdma_0_csr_write -> msgdma_0:csr_write
	wire   [31:0] mm_interconnect_1_msgdma_0_csr_writedata;                // mm_interconnect_1:msgdma_0_csr_writedata -> msgdma_0:csr_writedata
	wire          mm_interconnect_1_msgdma_0_descriptor_slave_waitrequest; // msgdma_0:descriptor_slave_waitrequest -> mm_interconnect_1:msgdma_0_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_1_msgdma_0_descriptor_slave_byteenable;  // mm_interconnect_1:msgdma_0_descriptor_slave_byteenable -> msgdma_0:descriptor_slave_byteenable
	wire          mm_interconnect_1_msgdma_0_descriptor_slave_write;       // mm_interconnect_1:msgdma_0_descriptor_slave_write -> msgdma_0:descriptor_slave_write
	wire  [127:0] mm_interconnect_1_msgdma_0_descriptor_slave_writedata;   // mm_interconnect_1:msgdma_0_descriptor_slave_writedata -> msgdma_0:descriptor_slave_writedata
	wire   [31:0] mm_interconnect_1_msgdma_0_response_readdata;            // msgdma_0:response_readdata -> mm_interconnect_1:msgdma_0_response_readdata
	wire          mm_interconnect_1_msgdma_0_response_waitrequest;         // msgdma_0:response_waitrequest -> mm_interconnect_1:msgdma_0_response_waitrequest
	wire    [0:0] mm_interconnect_1_msgdma_0_response_address;             // mm_interconnect_1:msgdma_0_response_address -> msgdma_0:response_address
	wire          mm_interconnect_1_msgdma_0_response_read;                // mm_interconnect_1:msgdma_0_response_read -> msgdma_0:response_read
	wire    [3:0] mm_interconnect_1_msgdma_0_response_byteenable;          // mm_interconnect_1:msgdma_0_response_byteenable -> msgdma_0:response_byteenable
	wire          msgdma_0_mm_write_waitrequest;                           // mm_interconnect_2:msgdma_0_mm_write_waitrequest -> msgdma_0:mm_write_waitrequest
	wire   [31:0] msgdma_0_mm_write_address;                               // msgdma_0:mm_write_address -> mm_interconnect_2:msgdma_0_mm_write_address
	wire    [7:0] msgdma_0_mm_write_byteenable;                            // msgdma_0:mm_write_byteenable -> mm_interconnect_2:msgdma_0_mm_write_byteenable
	wire          msgdma_0_mm_write_write;                                 // msgdma_0:mm_write_write -> mm_interconnect_2:msgdma_0_mm_write_write
	wire   [63:0] msgdma_0_mm_write_writedata;                             // msgdma_0:mm_write_writedata -> mm_interconnect_2:msgdma_0_mm_write_writedata
	wire          mm_interconnect_2_hps_0_f2h_sdram0_data_waitrequest;     // hps_0:f2h_sdram0_WAITREQUEST -> mm_interconnect_2:hps_0_f2h_sdram0_data_waitrequest
	wire   [28:0] mm_interconnect_2_hps_0_f2h_sdram0_data_address;         // mm_interconnect_2:hps_0_f2h_sdram0_data_address -> hps_0:f2h_sdram0_ADDRESS
	wire    [7:0] mm_interconnect_2_hps_0_f2h_sdram0_data_byteenable;      // mm_interconnect_2:hps_0_f2h_sdram0_data_byteenable -> hps_0:f2h_sdram0_BYTEENABLE
	wire          mm_interconnect_2_hps_0_f2h_sdram0_data_write;           // mm_interconnect_2:hps_0_f2h_sdram0_data_write -> hps_0:f2h_sdram0_WRITE
	wire   [63:0] mm_interconnect_2_hps_0_f2h_sdram0_data_writedata;       // mm_interconnect_2:hps_0_f2h_sdram0_data_writedata -> hps_0:f2h_sdram0_WRITEDATA
	wire    [7:0] mm_interconnect_2_hps_0_f2h_sdram0_data_burstcount;      // mm_interconnect_2:hps_0_f2h_sdram0_data_burstcount -> hps_0:f2h_sdram0_BURSTCOUNT
	wire          irq_mapper_receiver0_irq;                                // msgdma_0:csr_irq_irq -> irq_mapper:receiver0_irq
	wire   [31:0] hps_0_f2h_irq0_irq;                                      // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                      // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire          my_iq_source_0_avalon_streaming_source_valid;            // my_iq_source_0:stream_tvalid -> avalon_st_adapter:in_0_valid
	wire   [31:0] my_iq_source_0_avalon_streaming_source_data;             // my_iq_source_0:stream_tdata -> avalon_st_adapter:in_0_data
	wire          my_iq_source_0_avalon_streaming_source_ready;            // avalon_st_adapter:in_0_ready -> my_iq_source_0:stream_tready
	wire          my_iq_source_0_avalon_streaming_source_startofpacket;    // my_iq_source_0:stream_tstart -> avalon_st_adapter:in_0_startofpacket
	wire          my_iq_source_0_avalon_streaming_source_endofpacket;      // my_iq_source_0:stream_tlast -> avalon_st_adapter:in_0_endofpacket
	wire          avalon_st_adapter_out_0_valid;                           // avalon_st_adapter:out_0_valid -> dc_fifo_0:in_valid
	wire   [31:0] avalon_st_adapter_out_0_data;                            // avalon_st_adapter:out_0_data -> dc_fifo_0:in_data
	wire          avalon_st_adapter_out_0_ready;                           // dc_fifo_0:in_ready -> avalon_st_adapter:out_0_ready
	wire          avalon_st_adapter_out_0_startofpacket;                   // avalon_st_adapter:out_0_startofpacket -> dc_fifo_0:in_startofpacket
	wire          avalon_st_adapter_out_0_endofpacket;                     // avalon_st_adapter:out_0_endofpacket -> dc_fifo_0:in_endofpacket
	wire    [1:0] avalon_st_adapter_out_0_empty;                           // avalon_st_adapter:out_0_empty -> dc_fifo_0:in_empty
	wire          dc_fifo_0_out_valid;                                     // dc_fifo_0:out_valid -> avalon_st_adapter_001:in_0_valid
	wire   [31:0] dc_fifo_0_out_data;                                      // dc_fifo_0:out_data -> avalon_st_adapter_001:in_0_data
	wire          dc_fifo_0_out_ready;                                     // avalon_st_adapter_001:in_0_ready -> dc_fifo_0:out_ready
	wire          dc_fifo_0_out_startofpacket;                             // dc_fifo_0:out_startofpacket -> avalon_st_adapter_001:in_0_startofpacket
	wire          dc_fifo_0_out_endofpacket;                               // dc_fifo_0:out_endofpacket -> avalon_st_adapter_001:in_0_endofpacket
	wire    [1:0] dc_fifo_0_out_empty;                                     // dc_fifo_0:out_empty -> avalon_st_adapter_001:in_0_empty
	wire          avalon_st_adapter_001_out_0_valid;                       // avalon_st_adapter_001:out_0_valid -> msgdma_0:st_sink_valid
	wire   [63:0] avalon_st_adapter_001_out_0_data;                        // avalon_st_adapter_001:out_0_data -> msgdma_0:st_sink_data
	wire          avalon_st_adapter_001_out_0_ready;                       // msgdma_0:st_sink_ready -> avalon_st_adapter_001:out_0_ready
	wire          avalon_st_adapter_001_out_0_startofpacket;               // avalon_st_adapter_001:out_0_startofpacket -> msgdma_0:st_sink_startofpacket
	wire          avalon_st_adapter_001_out_0_endofpacket;                 // avalon_st_adapter_001:out_0_endofpacket -> msgdma_0:st_sink_endofpacket
	wire    [2:0] avalon_st_adapter_001_out_0_empty;                       // avalon_st_adapter_001:out_0_empty -> msgdma_0:st_sink_empty
	wire          rst_controller_reset_out_reset;                          // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, dc_fifo_0:in_reset_n, my_iq_source_0:reset]
	wire          rst_controller_001_reset_out_reset;                      // rst_controller_001:reset_out -> [avalon_st_adapter_001:in_rst_0_reset, dc_fifo_0:out_reset_n, mm_bridge_0:reset, mm_interconnect_0:mm_bridge_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:msgdma_0_reset_n_reset_bridge_in_reset_reset, mm_interconnect_2:msgdma_0_reset_n_reset_bridge_in_reset_reset, msgdma_0:reset_n_reset_n]
	wire          rst_controller_002_reset_out_reset;                      // rst_controller_002:reset_out -> [mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset]

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (4),
		.BITS_PER_SYMBOL    (8),
		.FIFO_DEPTH         (1024),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (1),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (3),
		.RD_SYNC_DEPTH      (3)
	) dc_fifo_0 (
		.in_clk            (lvds_clk_input_clk),                    //        in_clk.clk
		.in_reset_n        (~rst_controller_reset_out_reset),       //  in_clk_reset.reset_n
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset_n       (~rst_controller_001_reset_out_reset),   // out_clk_reset.reset_n
		.in_data           (avalon_st_adapter_out_0_data),          //            in.data
		.in_valid          (avalon_st_adapter_out_0_valid),         //              .valid
		.in_ready          (avalon_st_adapter_out_0_ready),         //              .ready
		.in_startofpacket  (avalon_st_adapter_out_0_startofpacket), //              .startofpacket
		.in_endofpacket    (avalon_st_adapter_out_0_endofpacket),   //              .endofpacket
		.in_empty          (avalon_st_adapter_out_0_empty),         //              .empty
		.out_data          (dc_fifo_0_out_data),                    //           out.data
		.out_valid         (dc_fifo_0_out_valid),                   //              .valid
		.out_ready         (dc_fifo_0_out_ready),                   //              .ready
		.out_startofpacket (dc_fifo_0_out_startofpacket),           //              .startofpacket
		.out_endofpacket   (dc_fifo_0_out_endofpacket),             //              .endofpacket
		.out_empty         (dc_fifo_0_out_empty),                   //              .empty
		.in_csr_address    (1'b0),                                  //   (terminated)
		.in_csr_read       (1'b0),                                  //   (terminated)
		.in_csr_write      (1'b0),                                  //   (terminated)
		.in_csr_readdata   (),                                      //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000),  //   (terminated)
		.out_csr_address   (1'b0),                                  //   (terminated)
		.out_csr_read      (1'b0),                                  //   (terminated)
		.out_csr_write     (1'b0),                                  //   (terminated)
		.out_csr_readdata  (),                                      //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000),  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_error         (),                                      //   (terminated)
		.in_channel        (1'b0),                                  //   (terminated)
		.out_channel       (),                                      //   (terminated)
		.space_avail_data  ()                                       //   (terminated)
	);

	soc_system_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.spim0_txd              (hps_0_spim0_f_txd),                                   //             spim0.txd
		.spim0_rxd              (hps_0_spim0_f_rxd),                                   //                  .rxd
		.spim0_ss_in_n          (hps_0_spim0_f_ss_in_n),                               //                  .ss_in_n
		.spim0_ssi_oe_n         (hps_0_spim0_f_ssi_oe_n),                              //                  .ssi_oe_n
		.spim0_ss_0_n           (hps_0_spim0_f_ss_0_n),                                //                  .ss_0_n
		.spim0_ss_1_n           (hps_0_spim0_f_ss_1_n),                                //                  .ss_1_n
		.spim0_ss_2_n           (hps_0_spim0_f_ss_2_n),                                //                  .ss_2_n
		.spim0_ss_3_n           (hps_0_spim0_f_ss_3_n),                                //                  .ss_3_n
		.spim0_sclk_out         (hps_0_spim0_sclk_out_f_clk),                          //    spim0_sclk_out.clk
		.mem_a                  (memory_mem_a),                                        //            memory.mem_a
		.mem_ba                 (memory_mem_ba),                                       //                  .mem_ba
		.mem_ck                 (memory_mem_ck),                                       //                  .mem_ck
		.mem_ck_n               (memory_mem_ck_n),                                     //                  .mem_ck_n
		.mem_cke                (memory_mem_cke),                                      //                  .mem_cke
		.mem_cs_n               (memory_mem_cs_n),                                     //                  .mem_cs_n
		.mem_ras_n              (memory_mem_ras_n),                                    //                  .mem_ras_n
		.mem_cas_n              (memory_mem_cas_n),                                    //                  .mem_cas_n
		.mem_we_n               (memory_mem_we_n),                                     //                  .mem_we_n
		.mem_reset_n            (memory_mem_reset_n),                                  //                  .mem_reset_n
		.mem_dq                 (memory_mem_dq),                                       //                  .mem_dq
		.mem_dqs                (memory_mem_dqs),                                      //                  .mem_dqs
		.mem_dqs_n              (memory_mem_dqs_n),                                    //                  .mem_dqs_n
		.mem_odt                (memory_mem_odt),                                      //                  .mem_odt
		.mem_dm                 (memory_mem_dm),                                       //                  .mem_dm
		.oct_rzqin              (memory_oct_rzqin),                                    //                  .oct_rzqin
		.h2f_rst_n              (hps_0_h2f_reset_reset_n),                             //         h2f_reset.reset_n
		.f2h_sdram0_clk         (clk_clk),                                             //  f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS     (mm_interconnect_2_hps_0_f2h_sdram0_data_address),     //   f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT  (mm_interconnect_2_hps_0_f2h_sdram0_data_burstcount),  //                  .burstcount
		.f2h_sdram0_WAITREQUEST (mm_interconnect_2_hps_0_f2h_sdram0_data_waitrequest), //                  .waitrequest
		.f2h_sdram0_WRITEDATA   (mm_interconnect_2_hps_0_f2h_sdram0_data_writedata),   //                  .writedata
		.f2h_sdram0_BYTEENABLE  (mm_interconnect_2_hps_0_f2h_sdram0_data_byteenable),  //                  .byteenable
		.f2h_sdram0_WRITE       (mm_interconnect_2_hps_0_f2h_sdram0_data_write),       //                  .write
		.h2f_axi_clk            (clk_clk),                                             //     h2f_axi_clock.clk
		.h2f_AWID               (hps_0_h2f_axi_master_awid),                           //    h2f_axi_master.awid
		.h2f_AWADDR             (hps_0_h2f_axi_master_awaddr),                         //                  .awaddr
		.h2f_AWLEN              (hps_0_h2f_axi_master_awlen),                          //                  .awlen
		.h2f_AWSIZE             (hps_0_h2f_axi_master_awsize),                         //                  .awsize
		.h2f_AWBURST            (hps_0_h2f_axi_master_awburst),                        //                  .awburst
		.h2f_AWLOCK             (hps_0_h2f_axi_master_awlock),                         //                  .awlock
		.h2f_AWCACHE            (hps_0_h2f_axi_master_awcache),                        //                  .awcache
		.h2f_AWPROT             (hps_0_h2f_axi_master_awprot),                         //                  .awprot
		.h2f_AWVALID            (hps_0_h2f_axi_master_awvalid),                        //                  .awvalid
		.h2f_AWREADY            (hps_0_h2f_axi_master_awready),                        //                  .awready
		.h2f_WID                (hps_0_h2f_axi_master_wid),                            //                  .wid
		.h2f_WDATA              (hps_0_h2f_axi_master_wdata),                          //                  .wdata
		.h2f_WSTRB              (hps_0_h2f_axi_master_wstrb),                          //                  .wstrb
		.h2f_WLAST              (hps_0_h2f_axi_master_wlast),                          //                  .wlast
		.h2f_WVALID             (hps_0_h2f_axi_master_wvalid),                         //                  .wvalid
		.h2f_WREADY             (hps_0_h2f_axi_master_wready),                         //                  .wready
		.h2f_BID                (hps_0_h2f_axi_master_bid),                            //                  .bid
		.h2f_BRESP              (hps_0_h2f_axi_master_bresp),                          //                  .bresp
		.h2f_BVALID             (hps_0_h2f_axi_master_bvalid),                         //                  .bvalid
		.h2f_BREADY             (hps_0_h2f_axi_master_bready),                         //                  .bready
		.h2f_ARID               (hps_0_h2f_axi_master_arid),                           //                  .arid
		.h2f_ARADDR             (hps_0_h2f_axi_master_araddr),                         //                  .araddr
		.h2f_ARLEN              (hps_0_h2f_axi_master_arlen),                          //                  .arlen
		.h2f_ARSIZE             (hps_0_h2f_axi_master_arsize),                         //                  .arsize
		.h2f_ARBURST            (hps_0_h2f_axi_master_arburst),                        //                  .arburst
		.h2f_ARLOCK             (hps_0_h2f_axi_master_arlock),                         //                  .arlock
		.h2f_ARCACHE            (hps_0_h2f_axi_master_arcache),                        //                  .arcache
		.h2f_ARPROT             (hps_0_h2f_axi_master_arprot),                         //                  .arprot
		.h2f_ARVALID            (hps_0_h2f_axi_master_arvalid),                        //                  .arvalid
		.h2f_ARREADY            (hps_0_h2f_axi_master_arready),                        //                  .arready
		.h2f_RID                (hps_0_h2f_axi_master_rid),                            //                  .rid
		.h2f_RDATA              (hps_0_h2f_axi_master_rdata),                          //                  .rdata
		.h2f_RRESP              (hps_0_h2f_axi_master_rresp),                          //                  .rresp
		.h2f_RLAST              (hps_0_h2f_axi_master_rlast),                          //                  .rlast
		.h2f_RVALID             (hps_0_h2f_axi_master_rvalid),                         //                  .rvalid
		.h2f_RREADY             (hps_0_h2f_axi_master_rready),                         //                  .rready
		.f2h_axi_clk            (clk_clk),                                             //     f2h_axi_clock.clk
		.f2h_AWID               (),                                                    //     f2h_axi_slave.awid
		.f2h_AWADDR             (),                                                    //                  .awaddr
		.f2h_AWLEN              (),                                                    //                  .awlen
		.f2h_AWSIZE             (),                                                    //                  .awsize
		.f2h_AWBURST            (),                                                    //                  .awburst
		.f2h_AWLOCK             (),                                                    //                  .awlock
		.f2h_AWCACHE            (),                                                    //                  .awcache
		.f2h_AWPROT             (),                                                    //                  .awprot
		.f2h_AWVALID            (),                                                    //                  .awvalid
		.f2h_AWREADY            (),                                                    //                  .awready
		.f2h_AWUSER             (),                                                    //                  .awuser
		.f2h_WID                (),                                                    //                  .wid
		.f2h_WDATA              (),                                                    //                  .wdata
		.f2h_WSTRB              (),                                                    //                  .wstrb
		.f2h_WLAST              (),                                                    //                  .wlast
		.f2h_WVALID             (),                                                    //                  .wvalid
		.f2h_WREADY             (),                                                    //                  .wready
		.f2h_BID                (),                                                    //                  .bid
		.f2h_BRESP              (),                                                    //                  .bresp
		.f2h_BVALID             (),                                                    //                  .bvalid
		.f2h_BREADY             (),                                                    //                  .bready
		.f2h_ARID               (),                                                    //                  .arid
		.f2h_ARADDR             (),                                                    //                  .araddr
		.f2h_ARLEN              (),                                                    //                  .arlen
		.f2h_ARSIZE             (),                                                    //                  .arsize
		.f2h_ARBURST            (),                                                    //                  .arburst
		.f2h_ARLOCK             (),                                                    //                  .arlock
		.f2h_ARCACHE            (),                                                    //                  .arcache
		.f2h_ARPROT             (),                                                    //                  .arprot
		.f2h_ARVALID            (),                                                    //                  .arvalid
		.f2h_ARREADY            (),                                                    //                  .arready
		.f2h_ARUSER             (),                                                    //                  .aruser
		.f2h_RID                (),                                                    //                  .rid
		.f2h_RDATA              (),                                                    //                  .rdata
		.f2h_RRESP              (),                                                    //                  .rresp
		.f2h_RLAST              (),                                                    //                  .rlast
		.f2h_RVALID             (),                                                    //                  .rvalid
		.f2h_RREADY             (),                                                    //                  .rready
		.h2f_lw_axi_clk         (clk_clk),                                             //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID            (hps_0_h2f_lw_axi_master_awid),                        // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR          (hps_0_h2f_lw_axi_master_awaddr),                      //                  .awaddr
		.h2f_lw_AWLEN           (hps_0_h2f_lw_axi_master_awlen),                       //                  .awlen
		.h2f_lw_AWSIZE          (hps_0_h2f_lw_axi_master_awsize),                      //                  .awsize
		.h2f_lw_AWBURST         (hps_0_h2f_lw_axi_master_awburst),                     //                  .awburst
		.h2f_lw_AWLOCK          (hps_0_h2f_lw_axi_master_awlock),                      //                  .awlock
		.h2f_lw_AWCACHE         (hps_0_h2f_lw_axi_master_awcache),                     //                  .awcache
		.h2f_lw_AWPROT          (hps_0_h2f_lw_axi_master_awprot),                      //                  .awprot
		.h2f_lw_AWVALID         (hps_0_h2f_lw_axi_master_awvalid),                     //                  .awvalid
		.h2f_lw_AWREADY         (hps_0_h2f_lw_axi_master_awready),                     //                  .awready
		.h2f_lw_WID             (hps_0_h2f_lw_axi_master_wid),                         //                  .wid
		.h2f_lw_WDATA           (hps_0_h2f_lw_axi_master_wdata),                       //                  .wdata
		.h2f_lw_WSTRB           (hps_0_h2f_lw_axi_master_wstrb),                       //                  .wstrb
		.h2f_lw_WLAST           (hps_0_h2f_lw_axi_master_wlast),                       //                  .wlast
		.h2f_lw_WVALID          (hps_0_h2f_lw_axi_master_wvalid),                      //                  .wvalid
		.h2f_lw_WREADY          (hps_0_h2f_lw_axi_master_wready),                      //                  .wready
		.h2f_lw_BID             (hps_0_h2f_lw_axi_master_bid),                         //                  .bid
		.h2f_lw_BRESP           (hps_0_h2f_lw_axi_master_bresp),                       //                  .bresp
		.h2f_lw_BVALID          (hps_0_h2f_lw_axi_master_bvalid),                      //                  .bvalid
		.h2f_lw_BREADY          (hps_0_h2f_lw_axi_master_bready),                      //                  .bready
		.h2f_lw_ARID            (hps_0_h2f_lw_axi_master_arid),                        //                  .arid
		.h2f_lw_ARADDR          (hps_0_h2f_lw_axi_master_araddr),                      //                  .araddr
		.h2f_lw_ARLEN           (hps_0_h2f_lw_axi_master_arlen),                       //                  .arlen
		.h2f_lw_ARSIZE          (hps_0_h2f_lw_axi_master_arsize),                      //                  .arsize
		.h2f_lw_ARBURST         (hps_0_h2f_lw_axi_master_arburst),                     //                  .arburst
		.h2f_lw_ARLOCK          (hps_0_h2f_lw_axi_master_arlock),                      //                  .arlock
		.h2f_lw_ARCACHE         (hps_0_h2f_lw_axi_master_arcache),                     //                  .arcache
		.h2f_lw_ARPROT          (hps_0_h2f_lw_axi_master_arprot),                      //                  .arprot
		.h2f_lw_ARVALID         (hps_0_h2f_lw_axi_master_arvalid),                     //                  .arvalid
		.h2f_lw_ARREADY         (hps_0_h2f_lw_axi_master_arready),                     //                  .arready
		.h2f_lw_RID             (hps_0_h2f_lw_axi_master_rid),                         //                  .rid
		.h2f_lw_RDATA           (hps_0_h2f_lw_axi_master_rdata),                       //                  .rdata
		.h2f_lw_RRESP           (hps_0_h2f_lw_axi_master_rresp),                       //                  .rresp
		.h2f_lw_RLAST           (hps_0_h2f_lw_axi_master_rlast),                       //                  .rlast
		.h2f_lw_RVALID          (hps_0_h2f_lw_axi_master_rvalid),                      //                  .rvalid
		.h2f_lw_RREADY          (hps_0_h2f_lw_axi_master_rready),                      //                  .rready
		.f2h_irq_p0             (hps_0_f2h_irq0_irq),                                  //          f2h_irq0.irq
		.f2h_irq_p1             (hps_0_f2h_irq1_irq)                                   //          f2h_irq1.irq
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (64),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (10),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (clk_clk),                                        //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),             // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (),                                               //    m0.waitrequest
		.m0_readdata      (),                                               //      .readdata
		.m0_readdatavalid (),                                               //      .readdatavalid
		.m0_burstcount    (),                                               //      .burstcount
		.m0_writedata     (),                                               //      .writedata
		.m0_address       (),                                               //      .address
		.m0_write         (),                                               //      .write
		.m0_read          (),                                               //      .read
		.m0_byteenable    (),                                               //      .byteenable
		.m0_debugaccess   (),                                               //      .debugaccess
		.s0_response      (),                                               // (terminated)
		.m0_response      (2'b00)                                           // (terminated)
	);

	soc_system_msgdma_0 msgdma_0 (
		.mm_write_address             (msgdma_0_mm_write_address),                               //         mm_write.address
		.mm_write_write               (msgdma_0_mm_write_write),                                 //                 .write
		.mm_write_byteenable          (msgdma_0_mm_write_byteenable),                            //                 .byteenable
		.mm_write_writedata           (msgdma_0_mm_write_writedata),                             //                 .writedata
		.mm_write_waitrequest         (msgdma_0_mm_write_waitrequest),                           //                 .waitrequest
		.clock_clk                    (clk_clk),                                                 //            clock.clk
		.reset_n_reset_n              (~rst_controller_001_reset_out_reset),                     //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_1_msgdma_0_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_1_msgdma_0_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_1_msgdma_0_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_1_msgdma_0_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_1_msgdma_0_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_1_msgdma_0_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_1_msgdma_0_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_1_msgdma_0_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_1_msgdma_0_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_1_msgdma_0_descriptor_slave_byteenable),  //                 .byteenable
		.response_waitrequest         (mm_interconnect_1_msgdma_0_response_waitrequest),         //         response.waitrequest
		.response_byteenable          (mm_interconnect_1_msgdma_0_response_byteenable),          //                 .byteenable
		.response_address             (mm_interconnect_1_msgdma_0_response_address),             //                 .address
		.response_readdata            (mm_interconnect_1_msgdma_0_response_readdata),            //                 .readdata
		.response_read                (mm_interconnect_1_msgdma_0_response_read),                //                 .read
		.csr_irq_irq                  (irq_mapper_receiver0_irq),                                //          csr_irq.irq
		.st_sink_data                 (avalon_st_adapter_001_out_0_data),                        //          st_sink.data
		.st_sink_valid                (avalon_st_adapter_001_out_0_valid),                       //                 .valid
		.st_sink_ready                (avalon_st_adapter_001_out_0_ready),                       //                 .ready
		.st_sink_startofpacket        (avalon_st_adapter_001_out_0_startofpacket),               //                 .startofpacket
		.st_sink_endofpacket          (avalon_st_adapter_001_out_0_endofpacket),                 //                 .endofpacket
		.st_sink_empty                (avalon_st_adapter_001_out_0_empty)                        //                 .empty
	);

	iq_stream_source_change #(
		.DATA_W (32)
	) my_iq_source_0 (
		.clk           (lvds_clk_input_clk),                                   //                   clock.clk
		.reset         (rst_controller_reset_out_reset),                       //                   reset.reset
		.stream_tdata  (my_iq_source_0_avalon_streaming_source_data),          // avalon_streaming_source.data
		.stream_tvalid (my_iq_source_0_avalon_streaming_source_valid),         //                        .valid
		.stream_tready (my_iq_source_0_avalon_streaming_source_ready),         //                        .ready
		.stream_tstart (my_iq_source_0_avalon_streaming_source_startofpacket), //                        .startofpacket
		.stream_tlast  (my_iq_source_0_avalon_streaming_source_endofpacket),   //                        .endofpacket
		.iq_word_in    (lvds_iq_hps_in_new_signal),                            //             conduit_end.new_signal
		.word_valid_in (word_valid_word_valid)                                 //           conduit_end_1.word_valid
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                      //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                    //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                     //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                    //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                   //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                    //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                   //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                    //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                   //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                   //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                       //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                     //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                     //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                     //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                    //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                    //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                       //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                     //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                    //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                    //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                      //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                    //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                     //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                    //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                   //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                    //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                   //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                    //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                   //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                   //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                       //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                     //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                     //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                     //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                    //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                    //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                        //                                                  clk_0_clk.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),             // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_reset_reset_bridge_in_reset_reset                    (rst_controller_001_reset_out_reset),             //                    mm_bridge_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_s0_address                                           (mm_interconnect_0_mm_bridge_0_s0_address),       //                                             mm_bridge_0_s0.address
		.mm_bridge_0_s0_write                                             (mm_interconnect_0_mm_bridge_0_s0_write),         //                                                           .write
		.mm_bridge_0_s0_read                                              (mm_interconnect_0_mm_bridge_0_s0_read),          //                                                           .read
		.mm_bridge_0_s0_readdata                                          (mm_interconnect_0_mm_bridge_0_s0_readdata),      //                                                           .readdata
		.mm_bridge_0_s0_writedata                                         (mm_interconnect_0_mm_bridge_0_s0_writedata),     //                                                           .writedata
		.mm_bridge_0_s0_burstcount                                        (mm_interconnect_0_mm_bridge_0_s0_burstcount),    //                                                           .burstcount
		.mm_bridge_0_s0_byteenable                                        (mm_interconnect_0_mm_bridge_0_s0_byteenable),    //                                                           .byteenable
		.mm_bridge_0_s0_readdatavalid                                     (mm_interconnect_0_mm_bridge_0_s0_readdatavalid), //                                                           .readdatavalid
		.mm_bridge_0_s0_waitrequest                                       (mm_interconnect_0_mm_bridge_0_s0_waitrequest),   //                                                           .waitrequest
		.mm_bridge_0_s0_debugaccess                                       (mm_interconnect_0_mm_bridge_0_s0_debugaccess)    //                                                           .debugaccess
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                            //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                          //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                           //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                          //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                         //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                          //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                         //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                          //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                         //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                         //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                             //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                           //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                           //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                           //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                          //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                          //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                             //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                           //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                          //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                          //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                            //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                          //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                           //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                          //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                         //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                          //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                         //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                          //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                         //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                         //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                             //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                           //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                           //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                           //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                          //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                          //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                                 //                                                     clk_0_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                      // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.msgdma_0_reset_n_reset_bridge_in_reset_reset                        (rst_controller_001_reset_out_reset),                      //                        msgdma_0_reset_n_reset_bridge_in_reset.reset
		.msgdma_0_csr_address                                                (mm_interconnect_1_msgdma_0_csr_address),                  //                                                  msgdma_0_csr.address
		.msgdma_0_csr_write                                                  (mm_interconnect_1_msgdma_0_csr_write),                    //                                                              .write
		.msgdma_0_csr_read                                                   (mm_interconnect_1_msgdma_0_csr_read),                     //                                                              .read
		.msgdma_0_csr_readdata                                               (mm_interconnect_1_msgdma_0_csr_readdata),                 //                                                              .readdata
		.msgdma_0_csr_writedata                                              (mm_interconnect_1_msgdma_0_csr_writedata),                //                                                              .writedata
		.msgdma_0_csr_byteenable                                             (mm_interconnect_1_msgdma_0_csr_byteenable),               //                                                              .byteenable
		.msgdma_0_descriptor_slave_write                                     (mm_interconnect_1_msgdma_0_descriptor_slave_write),       //                                     msgdma_0_descriptor_slave.write
		.msgdma_0_descriptor_slave_writedata                                 (mm_interconnect_1_msgdma_0_descriptor_slave_writedata),   //                                                              .writedata
		.msgdma_0_descriptor_slave_byteenable                                (mm_interconnect_1_msgdma_0_descriptor_slave_byteenable),  //                                                              .byteenable
		.msgdma_0_descriptor_slave_waitrequest                               (mm_interconnect_1_msgdma_0_descriptor_slave_waitrequest), //                                                              .waitrequest
		.msgdma_0_response_address                                           (mm_interconnect_1_msgdma_0_response_address),             //                                             msgdma_0_response.address
		.msgdma_0_response_read                                              (mm_interconnect_1_msgdma_0_response_read),                //                                                              .read
		.msgdma_0_response_readdata                                          (mm_interconnect_1_msgdma_0_response_readdata),            //                                                              .readdata
		.msgdma_0_response_byteenable                                        (mm_interconnect_1_msgdma_0_response_byteenable),          //                                                              .byteenable
		.msgdma_0_response_waitrequest                                       (mm_interconnect_1_msgdma_0_response_waitrequest)          //                                                              .waitrequest
	);

	soc_system_mm_interconnect_2 mm_interconnect_2 (
		.clk_0_clk_clk                                                      (clk_clk),                                             //                                                    clk_0_clk.clk
		.hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                  // hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
		.msgdma_0_reset_n_reset_bridge_in_reset_reset                       (rst_controller_001_reset_out_reset),                  //                       msgdma_0_reset_n_reset_bridge_in_reset.reset
		.msgdma_0_mm_write_address                                          (msgdma_0_mm_write_address),                           //                                            msgdma_0_mm_write.address
		.msgdma_0_mm_write_waitrequest                                      (msgdma_0_mm_write_waitrequest),                       //                                                             .waitrequest
		.msgdma_0_mm_write_byteenable                                       (msgdma_0_mm_write_byteenable),                        //                                                             .byteenable
		.msgdma_0_mm_write_write                                            (msgdma_0_mm_write_write),                             //                                                             .write
		.msgdma_0_mm_write_writedata                                        (msgdma_0_mm_write_writedata),                         //                                                             .writedata
		.hps_0_f2h_sdram0_data_address                                      (mm_interconnect_2_hps_0_f2h_sdram0_data_address),     //                                        hps_0_f2h_sdram0_data.address
		.hps_0_f2h_sdram0_data_write                                        (mm_interconnect_2_hps_0_f2h_sdram0_data_write),       //                                                             .write
		.hps_0_f2h_sdram0_data_writedata                                    (mm_interconnect_2_hps_0_f2h_sdram0_data_writedata),   //                                                             .writedata
		.hps_0_f2h_sdram0_data_burstcount                                   (mm_interconnect_2_hps_0_f2h_sdram0_data_burstcount),  //                                                             .burstcount
		.hps_0_f2h_sdram0_data_byteenable                                   (mm_interconnect_2_hps_0_f2h_sdram0_data_byteenable),  //                                                             .byteenable
		.hps_0_f2h_sdram0_data_waitrequest                                  (mm_interconnect_2_hps_0_f2h_sdram0_data_waitrequest)  //                                                             .waitrequest
	);

	soc_system_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	soc_system_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	soc_system_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (lvds_clk_input_clk),                                   // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),                       // in_rst_0.reset
		.in_0_data           (my_iq_source_0_avalon_streaming_source_data),          //     in_0.data
		.in_0_valid          (my_iq_source_0_avalon_streaming_source_valid),         //         .valid
		.in_0_ready          (my_iq_source_0_avalon_streaming_source_ready),         //         .ready
		.in_0_startofpacket  (my_iq_source_0_avalon_streaming_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (my_iq_source_0_avalon_streaming_source_endofpacket),   //         .endofpacket
		.out_0_data          (avalon_st_adapter_out_0_data),                         //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                        //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                        //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),                //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),                  //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty)                         //         .empty
	);

	soc_system_avalon_st_adapter_001 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (clk_clk),                                   // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_001_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (dc_fifo_0_out_data),                        //     in_0.data
		.in_0_valid          (dc_fifo_0_out_valid),                       //         .valid
		.in_0_ready          (dc_fifo_0_out_ready),                       //         .ready
		.in_0_startofpacket  (dc_fifo_0_out_startofpacket),               //         .startofpacket
		.in_0_endofpacket    (dc_fifo_0_out_endofpacket),                 //         .endofpacket
		.in_0_empty          (dc_fifo_0_out_empty),                       //         .empty
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_001_out_0_empty)          //         .empty
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (lvds_clk_input_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
