
module clkbuffer (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
